----------------------------------------------------------------------------------
-- Company: 
-- Engineer: Dordije Boskovic
-- 
-- Create Date: 
-- Design Name: 
-- Module Name: BRAM WRAPPER - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: Wrapper in VHDL because Vivado does not support VHDL 2008 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;

entity BRAM_WRAPPER is
	generic (

		-- Parameters of Axi Slave Bus Interface S00_AXI
		C_S00_AXI_DATA_WIDTH : integer := 25;
		C_S00_AXI_ADDR_WIDTH : integer := 4;

		--BRAM PARAMETERS
		BRAM_DATA_WIDTH      : integer := 25;
		NUM_BANDS            : integer := 16;
		BRAM_ADDR_WIDTH      : integer := 4 --integer(ceil(log2(real(NUM_BANDS))))
	);
	port (
		-- Users to add ports here

		-- User ports ends
		-- Do not modify the ports beyond this line
		-- Ports of Axi Slave Bus Interface S00_AXI
		s00_axi_aclk     : in std_logic;
		s00_axi_aresetn  : in std_logic;
		s00_axi_awaddr   : in std_logic_vector(C_S00_AXI_ADDR_WIDTH - 1 downto 0);
		s00_axi_awprot   : in std_logic_vector(2 downto 0);
		s00_axi_awvalid  : in std_logic;
		s00_axi_awready  : out std_logic;
		s00_axi_wdata    : in std_logic_vector(C_S00_AXI_DATA_WIDTH - 1 downto 0);
		s00_axi_wstrb    : in std_logic_vector((C_S00_AXI_DATA_WIDTH/8) - 1 downto 0);
		s00_axi_wvalid   : in std_logic;
		s00_axi_wready   : out std_logic;
		s00_axi_bresp    : out std_logic_vector(1 downto 0);
		s00_axi_bvalid   : out std_logic;
		s00_axi_bready   : in std_logic;
		s00_axi_araddr   : in std_logic_vector(C_S00_AXI_ADDR_WIDTH - 1 downto 0);
		s00_axi_arprot   : in std_logic_vector(2 downto 0);
		s00_axi_arvalid  : in std_logic;
		s00_axi_arready  : out std_logic;
		s00_axi_rdata    : out std_logic_vector(C_S00_AXI_DATA_WIDTH - 1 downto 0);
		s00_axi_rresp    : out std_logic_vector(1 downto 0);
		s00_axi_rvalid   : out std_logic;
		s00_axi_rready   : in std_logic;

		--BRAM SIGNALS
		MATRIX_ROW       : out std_logic_vector(BRAM_DATA_WIDTH * NUM_BANDS - 1 downto 0);
		ROW_SELECT       : in std_logic_vector (BRAM_ADDR_WIDTH - 1 downto 0);
		STATIC_VECTOR_SR : out std_logic_vector (BRAM_DATA_WIDTH - 1 downto 0)
	);
end BRAM_WRAPPER;

architecture arch_imp of BRAM_WRAPPER is

	-- component declaration
	component AXI_BRAM is
		generic (
			C_S_AXI_DATA_WIDTH : integer := 32;
			-- Width of S_AXI address bus
			C_S_AXI_ADDR_WIDTH : integer := 4;
			--BRAM PARAMETERS
			BRAM_DATA_WIDTH    : integer := 32;
			NUM_BANDS          : integer := 16;
			BRAM_ADDR_WIDTH    : integer := 4--integer(ceil(log2(real(NUM_BANDS))))
		);
		port (
			S_AXI_ACLK       : in std_logic;
			S_AXI_ARESETN    : in std_logic;
			S_AXI_AWADDR     : in std_logic_vector(C_S_AXI_ADDR_WIDTH - 1 downto 0);
			S_AXI_AWPROT     : in std_logic_vector(2 downto 0);
			S_AXI_AWVALID    : in std_logic;
			S_AXI_AWREADY    : out std_logic;
			S_AXI_WDATA      : in std_logic_vector(C_S_AXI_DATA_WIDTH - 1 downto 0);
			S_AXI_WSTRB      : in std_logic_vector((C_S_AXI_DATA_WIDTH/8) - 1 downto 0);
			S_AXI_WVALID     : in std_logic;
			S_AXI_WREADY     : out std_logic;
			S_AXI_BRESP      : out std_logic_vector(1 downto 0);
			S_AXI_BVALID     : out std_logic;
			S_AXI_BREADY     : in std_logic;
			S_AXI_ARADDR     : in std_logic_vector(C_S_AXI_ADDR_WIDTH - 1 downto 0);
			S_AXI_ARPROT     : in std_logic_vector(2 downto 0);
			S_AXI_ARVALID    : in std_logic;
			S_AXI_ARREADY    : out std_logic;
			S_AXI_RDATA      : out std_logic_vector(C_S_AXI_DATA_WIDTH - 1 downto 0);
			S_AXI_RRESP      : out std_logic_vector(1 downto 0);
			S_AXI_RVALID     : out std_logic;
			S_AXI_RREADY     : in std_logic;
			MATRIX_ROW       : out std_logic_vector(BRAM_DATA_WIDTH * NUM_BANDS - 1 downto 0);
			ROW_SELECT       : in std_logic_vector (BRAM_ADDR_WIDTH - 1 downto 0);
			STATIC_VECTOR_SR : out std_logic_vector (BRAM_DATA_WIDTH - 1 downto 0)
		);
	end component AXI_BRAM;

begin

	-- Instantiation of Axi Bus Interface S00_AXI
	AXI_BRAM_inst : AXI_BRAM
	generic map(
		C_S_AXI_DATA_WIDTH => C_S00_AXI_DATA_WIDTH,
		C_S_AXI_ADDR_WIDTH => C_S00_AXI_ADDR_WIDTH,
		BRAM_DATA_WIDTH    => BRAM_DATA_WIDTH,
		NUM_BANDS          => NUM_BANDS,
		BRAM_ADDR_WIDTH    => BRAM_ADDR_WIDTH
	)
	port map(
		S_AXI_ACLK       => s00_axi_aclk,
		S_AXI_ARESETN    => s00_axi_aresetn,
		S_AXI_AWADDR     => s00_axi_awaddr,
		S_AXI_AWPROT     => s00_axi_awprot,
		S_AXI_AWVALID    => s00_axi_awvalid,
		S_AXI_AWREADY    => s00_axi_awready,
		S_AXI_WDATA      => s00_axi_wdata,
		S_AXI_WSTRB      => s00_axi_wstrb,
		S_AXI_WVALID     => s00_axi_wvalid,
		S_AXI_WREADY     => s00_axi_wready,
		S_AXI_BRESP      => s00_axi_bresp,
		S_AXI_BVALID     => s00_axi_bvalid,
		S_AXI_BREADY     => s00_axi_bready,
		S_AXI_ARADDR     => s00_axi_araddr,
		S_AXI_ARPROT     => s00_axi_arprot,
		S_AXI_ARVALID    => s00_axi_arvalid,
		S_AXI_ARREADY    => s00_axi_arready,
		S_AXI_RDATA      => s00_axi_rdata,
		S_AXI_RRESP      => s00_axi_rresp,
		S_AXI_RVALID     => s00_axi_rvalid,
		S_AXI_RREADY     => s00_axi_rready,
		MATRIX_ROW       => MATRIX_ROW,
		ROW_SELECT       => ROW_SELECT,
		STATIC_VECTOR_SR => STATIC_VECTOR_SR
	);

	-- Add user logic here

	-- User logic ends

end arch_imp;